module memoria (clock, escrever, endereco, din, dout);

  input clock, escrever;
  input [15:0] endereco, din;
  output [15:0] dout;

  reg [15:0] mem [0:63]; // 64 x 16

  initial begin
    // Teste 1
    mem[0] <= 16'b1001100000000000;     // MVI  R4 #38
    mem[1] <= 16'b0000000000100110;     // #38
    mem[2] <= 16'b1001000000000000;     // MVI  R0 #2
    mem[3] <= 16'b0000000000000010;     // #2
    mem[4] <= 16'b1001001000000000;     // MVI  R1 #3
    mem[5] <= 16'b0000000000000011;     // #3
    mem[6] <= 16'b0000001000000000;     // ADD  R1 R0
    mem[7] <= 16'b1001010000000000;     // MVI  R2 #6
    mem[8] <= 16'b0000000000000110;     // #6
    mem[9] <= 16'b0001010001000000;     // SUB  R2 R1
    mem[10] <= 16'b1000011010000000;    // MV   R3 R2
    mem[11] <= 16'b0000000011000000;    // ADD  R0 R3
    mem[12] <= 16'b0010000001000000;    // AND  R0 R1
    mem[13] <= 16'b0100001011000000;    // SLL  R1 R3
    mem[14] <= 16'b0101001011000000;    // SRL  R1 R3
    mem[15] <= 16'b1001000000000000;    // MVI  R0 #0
    mem[16] <= 16'b0000000000000000;    // #0
    mem[17] <= 16'b0011000001000000;    // SLT  R0 R1
    mem[18] <= 16'b0011001001000000;    // SLT  R1 R1
    mem[19] <= 16'b1001011000000000;    // MVI  R3 #3
    mem[20] <= 16'b0000000000000011;    // #3
    mem[21] <= 16'b1001001000000000;    // MVI  R1 #5
    mem[22] <= 16'b0000000000000101;    // #5
    mem[23] <= 16'b0000000011000000;    // ADD  R0 R3
    mem[24] <= 16'b1001000000000000;    // MVI  R0 #0
    mem[25] <= 16'b0000000000000000;    // #0
    mem[26] <= 16'b0111010100000000;    // LD   R2 R4                 ** comando modificado **
    mem[27] <= 16'b0000010011000000;    // ADD  R2 R3
    mem[28] <= 16'b0110010000000000;    // SD   R2 R0
    mem[29] <= 16'b0111000000000000;    // LD   R0 R0
    mem[30] <= 16'b0001000011000000;    // SUB  R0 R3
    mem[31] <= 16'b1001000000000000;    // MVI  R0 #0
    mem[32] <= 16'b0000000000000000;    // #0
    mem[33] <= 16'b0000000000000000;    // ADD  R0 R0
    mem[34] <= 16'b1010000010000000;    // MVNZ R0 R2
    mem[35] <= 16'b0001001011000000;    // SUB  R1 R3
    mem[36] <= 16'b1010000010000000;    // MVNZ R0 R2
    mem[37] <= 16'b0000000001000000;    // ADD  R0 R1
    mem[38] <= 16'b0000000000000100;    // #4

    /*
    // Teste 2
    mem[0] <= 16'b1001010000000000;
    mem[1] <= 16'b0000000000000001;
    mem[2] <= 16'b1001100000000000;
    mem[3] <= 16'b0000000000001010;
    mem[4] <= 16'b1000101111000000;
    mem[5] <= 16'b0001100010000000;
    mem[6] <= 16'b1010111101000000;
    */
  end

  // Sempre realiza a leitura (assincrona)
  assign dout = mem[endereco];

  always @(posedge clock)
    if(escrever)
      mem[endereco] <= din;

endmodule
